
module ALU(input reg opcode, operand1, operand2, statusIn 
           output reg result, statusOut);
   
endmodule; // ALU

module testbench();
   
endmodule; // testbench

